Test Prob in class

v1 1 2 1
v2 3 0 2
v3 4 3 3

i1 0 3 1

r2 2 3 1
r1 1 0 1
r3 3 4 1
r4 0 3 1
r5 5 4 1 

.op
.tran 1us 100us
.control
run
write 
display 
print all
.endc

.end
