***Audio Ampilfier***

Vin 0 1 dc 0V ac sin(0 1 1kHz)
V1 8 0  dc 12V
V2 0 6 dc 12V

R4 2 0 100k
R5 7 3 510
R1 4 5 1k
R3 5 6 6.5k
R6 8 7 1k
R2 9 5 1k
R7 8 10 1.5k
R8 13 16 10k
R9 13 12 100k
R11 14 6 1k
R12 18 12 1
R13 12 0 8
R10 12 15 1

C1 1 2 2.2u
C2 16 0 47u

D1 11 17 D1N4500
D2 17 19 D1N4500
D3 19 14 D1N4500

Q1 3 2 4 Q2N3904
Q2 10 13 9 Q2N3904
Q3 11 7 8 Q2N3906
Q4 8 11 18 Qtip29
Q5 6 14 15 Qtip30 

.SUBCKT D1N4500 1 2
D1	1	2	DFWD
D1A	1	2	DXTRA
D1B	2	1	DLEAK
R	1	2	1.66407G

.MODEL DFWD D(IS=71.94942E-15 N=0.960183 RS=0.236317 IKF=0.000237528 CJO=4.0000E-12 M=.3333 VJ=.75 ISR=96.49884E-15 NR=1.82557 BV=86.542 IBV=.3447 TT=6.6562E-9)

.MODEL DXTRA D(IS = 68.81973E-12 RS = 28.47153E-3 N = 2.15458 IKF = 0.0531356 TT = 0 CJO = 0 VJ = 1 M = .5 EG = 1.11 XTI = 3 KF = 0 AF = 1 FC = .5 BV = 1E5 IBV = .001)

.MODEL DLEAK D(IS = 5.810722E-15 RS = 0.1 N = 180.584 TT = 0 CJO = 0 VJ = 1 M = .5 EG = 1.11 XTI = 3 KF = 0 AF = 1 FC = .5 BV = 1E5 IBV = .001
.ENDS
     
.MODEL Q2N3904	NPN(Is=6.734f Xti=3 Eg=1.11 Vaf=74.03 Bf=416.4 Ne=1.259 Ise=6.734f Ikf=66.78m Xtb=1.5 Br=.7371 Nc=2 Isc=0 Ikr=0 Rc=1 Cjc=3.638p Mjc=.3085 Vjc=.75 Fc=.5 Cje=4.493p Mje=.2593 Vje=.75 Tr=239.5n Tf=301.2p Itf=.4 Vtf=4 Xtf=2 Rb=10)
.MODEL Q2N3906  PNP (IS=7.9190E-15 BF=196.89 VAF=100 IKF=.7271 ISE=13.654E-15 NE=1.4535 BR=124.61 VAR=100 IKR=10.010E-3 ISC=18.518E-12 NC=1.6031 NK=1.1475 RB=8.6624 RC=.55428 CJE=11.640E-12 VJE=1.0397 MJE=.47196 CJC=7.8722E-12 VJC=.98301 MJC=.53872 TF=320.13E-12 XTF=29.514 VTF=81.870 ITF=.12448 TR=10.000E-9)
.MODEL Qtip29 NPN(IS=1e-09 BF=331.58 NF=0.85 VAF=52.0929 IKF=0.286747 ISE=1.27813e-09 NE=1.29493 BR=1.03668 NR=0.75 VAR=91.9558 IKR=1.91753 ISC=1.27813e-09 NC=3.05613 RB=43.0821 IRB=0.1 RBM=0.122668 RE=0.000563203 RC=0.34452 XTB=0.720859 XTI=1.14559 EG=1.05 CJE=7.7589e-08 VJE=0.550883 MJE=0.500345 TF=1e-08 XTF=1.35725 VTF=0.996005 ITF=0.999927 CJC=4.44553e-10 VJC=0.400343 MJC=0.409703 XCJC=0.803124 FC=0.568788 CJS=0 VJS=0.75 MJS=0.5 TR=1e-07 PTF=0 KF=0 AF=1)
.MODEL Qtip30 PNP(IS=1e-09 BF=192.893 NF=0.85 VAF=49.329 IKF=0.519667 ISE=1e-08 NE=1.90927 BR=1.14712 NR=1.5 VAR=58.8376 IKR=5.19667 ISC=1e-08 NC=3.07207 RB=45.4356 IRB=0.1 RBM=0.115769 RE=0.000526622 RC=0.718902 XTB=0.771093 XTI=1.16111 EG=1.05 CJE=8.27904e-08 VJE=0.538348 MJE=0.517133 TF=1e-08 XTF=1.35724 VTF=0.995977 ITF=0.999928 CJC=4.44657e-10 VJC=0.400388 MJC=0.409559 XCJC=0.803124 FC=0.571623 CJS=0 VJS=0.75 MJS=0.5 TR=1e-07 PTF=0 KF=0 AF=1)


.tran 1us 10ms
.control
run
write
display
.endc
.end
